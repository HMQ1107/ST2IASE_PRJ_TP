module linear_reg (size,prize,cout);
    input [15:0] size;
    input [15:0] price;

    output [31:0] cout;


endmodule : linear_reg