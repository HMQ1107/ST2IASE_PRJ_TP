module multiplier_16bit (a,b,cout);
    input [15:0] a;
    input [15:0] b;

    output [31:0] cout;


endmodule : multiplier_16bit